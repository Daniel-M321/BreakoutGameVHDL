-- Description: breakout game component
-- FSM-based design 

-- Engineer: Fearghal Morgan, National University of Ireland, Galway
-- Date: 26/10/2022
-- 
-- 16 x 32-bit game array, using reg32x32(15 downto 0)(31:0)

-- On completion
--    write reg4x32_CSRA(0)(1:0)  = 0b10, i.e, (1) = 1 => FPGA done, (0) = 0 => return control to host. Other CSRA(0) bits unchanged
--
-- Signal dictionary
--  clk					system clock strobe, rising edge active
--  rst	        		assertion (h) asynchronously clears all registers
--  ce                  chip enable, asserted high                 		 
--  go			        Assertion (H) detected in idle state to active threshold function 
--  active (Output)     Default asserted (h), except in idle state

--  reg4x32_CSRA    	4 x 32-bit Control & Status registers, CSRA
--  reg4x32_CSRB      	32-bit Control register, CSRB
--  BRAM_dOut	        Current source memory 256-bit data (not used in this application)

--  wr  (Output)        Asserted to synchronously write to addressed memory
--  add (Output)  	    Addressed memory - 0b00100000 to read BRAM(255:0)
--  datToMem (Output)   32-bit data to addressed memory 

--  functBus            96-bit array of function signals, for use in debug and demonstration of function behaviour 
--  			        Not used in this example

-- Internal Signal dictionary
--  NS, CS                         finite state machine state signals 
--  NS*, CS* 				       next and current state signals 

--    Using integer types for INTERNAL address signals where possible, to make VHDL model more readable

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.arrayPackage.all;

entity game is
    Port ( clk 		     : in STD_LOGIC;   
           rst 		     : in STD_LOGIC; 
           ce            : in  std_logic;                		 
           go            : in  std_logic;                		 
		   active        : out std_logic;

		   reg4x32_CSRA  : in array4x32; 
		   reg4x32_CSRB  : in array4x32;	
           BRAM_dOut     : in std_logic_vector(255 downto 0);	
           reg32x32_dOut : in std_logic_vector(31 downto 0);
					 
		   wr            : out std_logic;
		   add           : out std_logic_vector(  7 downto 0);					 
		   datToMem	     : out std_logic_vector( 31 downto 0);

		   functBus      : out std_logic_vector(95 downto 0)
           );
end game;

architecture RTL of game is
-- Internal signal declarations
-- <include new states>
type stateType is (idle, writeToCSR0, setupGameParameters, initGameArena, initBall, initPaddle, initLives, initScore, waitState, processPaddle, processBall, writeBallToMem, writeWallToMem, endGame, NW, N, NE, SE, S, SW); -- declare enumerated state type
signal NS, CS                                   : stateType; -- declare FSM state 
								                
signal NSWallVec, CSWallVec                     : std_logic_vector(31 downto 0);
signal NSBallVec, CSBallVec                     : std_logic_vector(31 downto 0);
signal NSPaddleVec, CSPaddleVec                 : std_logic_vector(31 downto 0);
								                
signal NSBallXAdd, CSBallXAdd                   : integer range 0 to 31;
signal NSBallYAdd, CSBallYAdd                   : integer range 0 to 31;
signal NSBallDir, CSBallDir                     : std_logic_vector(2 downto 0);
								                
signal NSScore, CSScore                         : integer range 0 to 31;
signal NSLives, CSLives                         : integer range 0 to 31;

-- Clock frequency = 12.5MHz, count 0 - 12,499,999 to create 1 second delay 
-- 100ms delay => count ~ 0 - 1,250,000
signal NSDlyCountMax, CSDlyCountMax             : integer range 0 to 1250000;
signal NSDlyCount, CSDlyCount                   : integer range 0 to 1250000;

signal NSPaddleNumDlyMax, CSPaddleNumDlyMax     : integer range 0 to 31;
signal NSPaddleNumDlyCount, CSPaddleNumDlyCount : integer range 0 to 31;

signal NSBallNumDlyMax, CSBallNumDlyMax         : integer range 0 to 31;
signal NSBallNumDlyCount, CSBallNumDlyCount     : integer range 0 to 31;

signal zone 									: integer; 

begin

asgnFunctBus2_i: functBus <= (others => '0'); -- not currently used 

-- FSM next state and o/p decode process
-- <include new signals in sensitivity list>
NSAndOPDec_i: process (CS, go, 
					   reg4x32_CSRA, reg4x32_CSRB, reg32x32_dOut, 
					   CSWallVec, CSPaddleVec, CSBallXAdd, CSBallYAdd, CSBallDir, CSScore, CSLives, 
					   CSDlyCountMax, CSPaddleNumDlyMax, CSBallNumDlyMax, CSDlyCount, CSPaddleNumDlyCount, CSBallNumDlyCount)
begin
   NS 	 		       <= CS;     -- default signal assignments
   NSWallVec           <= CSWallVec;
   NSBallVec           <= CSBallVec;
   NSPaddleVec         <= CSPaddleVec;
   NSBallXAdd          <= CSBallXAdd;
   NSBallYAdd          <= CSBallYAdd;
   NSBallDir           <= CSBallDir;
   NSScore             <= CSScore;
   NSLives             <= CSLives;
   NSDlyCount          <= CSDlyCount;           
   NSPaddleNumDlyCount <= CSPaddleNumDlyCount;
   NSBallNumDlyCount   <= CSBallNumDlyCount; 
   NSDlyCountMax       <= CSDlyCountMax;
   NSDlyCount          <= CSDlyCount;
   NSPaddleNumDlyMax   <= CSPaddleNumDlyMax;
   NSBallNumDlyMax     <= CSBallNumDlyMax;
   active    	       <= '1';             -- default asserted. Deasserted only in idle state. 
   wr   	           <= '0';
   add	               <= "010" & "00000"; -- reg32x32 base address
   datToMem            <= (others => '0');
   zone                <= 0;

  case CS is 
		when idle => 			     
			active  <= '0';  
            if go = '1' then 
				if    reg4x32_CSRA(0)(10 downto 8) = "000" then -- initialise game values and progress to init game arena states 
					NS 					<= setupGameParameters;							
				elsif reg4x32_CSRA(0)(10 downto 8) = "001" then -- play game
					NSDlyCount          <= 0;                   -- clear delay counters  
					NSPaddleNumDlyCount <= 0;  
					NSBallNumDlyCount   <= 0;
					NS                  <= waitState;
				end if;
			end if;

		when writeToCSR0 =>                                        -- finish. Return done state and return control to host
			wr       <= '1';
            add      <= "000" & "00000"; 						   -- reg4x32_CSRA address = 0 
		    datToMem <=   reg4x32_CSRA(0)(31 downto  8)            -- bits unchanged 
                        & reg4x32_CSRA(0)( 7 downto  2) & "10";    -- byte 0, bit(1) = 1 => FPGA done, bit(0) = 0 => return control to host. Bits 7:2 unchanged
			NS       <= idle;


		when setupGameParameters =>  
			NSWallVec           <= reg4x32_CSRA(3);
			NSBallXAdd 	        <= to_integer( unsigned(reg4x32_CSRA(2)(28 downto 24)) );
			NSBallYAdd 	        <= to_integer( unsigned(reg4x32_CSRA(2)(20 downto 16)) );
			NSLives             <= to_integer( unsigned(reg4x32_CSRA(2)( 3 downto  0)) );
			NSScore             <= to_integer( unsigned(reg4x32_CSRA(2)( 7 downto  4)) );
			NSBallVec           <= reg4x32_CSRA(1);

			NSPaddleVec         <= reg4x32_CSRB(3);
			NSBallDir           <= reg4x32_CSRB(2)(26 downto  24);
			NSDlyCountMax       <= to_integer( unsigned(reg4x32_CSRB(2)(19 downto  0)) );                 
			NSPaddleNumDlyMax   <= to_integer( unsigned(reg4x32_CSRB(1)(28 downto 24)) );
			NSBallNumDlyMax     <= to_integer( unsigned(reg4x32_CSRB(1)(20 downto 16)) );
			NS                  <= initGameArena;

		when initGameArena => -- follow an initialisation sequence              TODO where do these initial values come from? Is wallVec actaully full of 1s?
            -- write wallVec
			wr   	      <= '1';
			add           <= "010" & "01111";               -- reg32x32 row 15
			datToMem      <= CSWallVec;
           	NS            <= initBall;
        when initLives =>                          
			wr   	      <= '1';
			add	          <= "010" & "00001";               -- reg32x32 row 1
			datToMem      <= X"000000" & "000" & std_logic_vector( to_unsigned(CSLives, 5) );  
           	NS            <= initScore;     
		when initScore =>                          
			wr   	      <= '1';
			add	          <= "010" & "00000";               -- reg32x32 row 0 
			datToMem      <= X"000000" & "000" & std_logic_vector( to_unsigned(CSScore, 5) );  
           	NS            <= initBall;
		when initBall =>                                                                              -- DAN switched these around for when reseting round
			wr   	      <= '1';
			add	          <= "010" & std_logic_vector( to_unsigned(CSBallYAdd,5) );  
			datToMem      <= CSBallVec;
           	NS            <= initPaddle;
		when initPaddle =>
			wr   	      <= '1';
			add	          <= "010" & "00010";               -- reg32x32 row 2 
			datToMem      <= CSPaddleVec;
           	NS            <= writeToCSR0;                   -- finish. Return done state and return control to host


		when waitState =>                                   -- increment count and loop in state until value reaches delay value       
			if CSDlyCount = CSDlyCountMax then
	     	    NSDlyCount <= 0;                            -- clear delay counter and process paddle and/or ball	     	         	    
   	   	        NS  <= processPaddle;
            else
	   	        NSDlyCount    <= CSDlyCount + 1;                
			end if;
			
	     	    			
        -- read reg4x32_CSRA(0)(9:8) and move paddle left / right, between boundaries
		when processPaddle =>                               -- read CSRB(0)(9:8)
			if CSPaddleNumDlyCount = CSPaddleNumDlyMax then
	     	   NSPaddleNumDlyCount <= 0;                    -- clear counter
		       add	<= "010" & "00010";                     -- reg32x32 row 2 (paddle row) 
			     if reg4x32_CSRB(0)(9) = '1' then           -- if 1 in (9) -> shift paddle left, if not at bit 31 boundary
			        if reg32x32_dOut(31) = '0' then 
				        wr   	      <= '1';
					    add	          <= "010" & "00010";   -- reg32x32 row 2, paddle row address 
					    datToMem      <= reg32x32_dOut(30 downto 0) & '0'; 
				    end if;
			      elsif reg4x32_CSRB(0)(8) = '1' then       -- if 1 in (8) -> shift paddle right 
			        if reg32x32_dOut(0) = '0' then 
					    wr   	      <= '1';
					    add	          <= "010" & "00010";   -- reg32x32 row 2, paddle row address 
					    datToMem      <= '0' & reg32x32_dOut(31 downto 1); 
				    end if;
				  end if;   		  
           	else
	           NSPaddleNumDlyCount <= CSPaddleNumDlyCount + 1; -- increment counter
           	   NS  <= processBall;
           	end if;		

		-- ========= Only partially completed =========
        when processBall => 	
			if CSBallNumDlyCount = CSBallNumDlyMax then
		   	   NSBallNumDlyCount   <= 0;

               -- < instructions>		      
			   -- Perform ball zone checks with respect to boundaries, wall, paddle. 
			   -- Assign signal zone, for reference only
		       -- Update ball X/Y, directon, score, lives, wall. 
		       -- Check if end game
	 	       -- loop to waitState or progress to endGame
		
			   -- Check if ZoneCentral Y4To13_X1To30, up or down  
			   
			   -- Step 1 find the zone in this state, we have 
			   if CSBallYAdd >= 4 and CSBallYAdd <= 13 and CSBallXAdd >= 1 and CSBallXAdd <= 30 then  
			      zone <= 1;
				  if CSBallDir(2) = '1' then                        -- ball direction is up                               -- ball direction is up?
			         NSBallYAdd                  <= CSBallYAdd + 1; -- move up in Y direction
                     case CSBallDir(1 downto 0) is                                               -- 00 no CSBallXAdd change, 11 not valid, will not occur
                       when "01"   => NSBallXAdd <= CSBallXAdd - 1;                              -- if NE, decrement NSBallXAdd, moving east 
                       when "10"   => NSBallXAdd <= CSBallXAdd + 1;                              -- if NW, increment XAdd, moving west 
                       when others => null;                                                      -- no change
                     end case;                                                           
			       else  						                    -- ball direction is down                             -- ball direction is down?
			         NSBallYAdd                  <= CSBallYAdd - 1;                              -- move down in Y direction		 
                     case CSBallDir(1 downto 0) is                                               -- 00 no CSBallXAdd change, 11 not valid, will not occur
                       when "01"   => NSBallXAdd <= CSBallXAdd - 1;                              -- if SE, decrement NSBallXAdd, moving east 
                       when "10"   => NSBallXAdd <= CSBallXAdd + 1;                              -- if SW, increment NSBallXAdd, moving west 
                       when others => null; 									                 -- no change
                     end case;
			       end if;
                   wr                  <= '1'; 					        			             -- clear current ball row
                   add(7 downto 5)     <= "010";                                                 -- reg32x32 memory bank select 
                   add(4 downto 0)     <= std_logic_vector( to_unsigned(CSBallYAdd, 5) );        -- current row address 
	   		       datToMem            <= (others => '0');							             -- clear row
				   NS                  <= writeBallToMem;
			   
--			   elsif CSBallYAdd = 15 then                                                         -- zone 6, inside wall zone
--			       zone <= 6;
--			       if CSBallXAdd = 0 then
--			           NSBallXAdd <= CSBallXAdd + 1;
--			           NSBallYAdd <= CSBallYAdd - 1;
--			       elsif CSBallXAdd = 31 then
--			           NSBallXAdd <= CSBallXAdd - 1;
--			           NSBallYAdd <= CSBallYAdd - 1;
--			       if CSBallDir(2) = '1' then
--			           case CSBallDir(1 downto 0) is                                               -- 00 no CSBallXAdd change, 11 not valid, will not occur
--                         when "01"   => NSBallXAdd <= CSBallXAdd - 1;                              -- if NE, decrement NSBallXAdd, moving east 
--                         when "10"   => NSBallXAdd <= CSBallXAdd + 1;                              -- if NW, increment XAdd, moving west 
--                         when others => null;                                                      -- no change
--                       end case; 

               elsif CSBallXAdd = 31 then                                                       -- left wall
                   if CSBallYAdd = 4 then                                                       -- above paddle in left corner
                      zone <= 7;
                      add	<= "010" & "00010";                                                 -- paddle row
                      if reg32x32_dOut(31) = '1' then                                           -- if paddle
                          NSBallXAdd <= CSBallXAdd - 1;                                         -- NE
             	          NSBallYAdd <= CSBallYAdd + 1;
             	          NsBallDir <= "101";
             	      else                                                                      -- else lose a life
             	          NSLives <= CSLives - 1;
             	          if NSLives > 0 then                                                   -- TODO Is ballVec being updated anywhere?
             	              NS <= initBall;
             	              NSBallXAdd <= 16;                                                 -- ball back to middle above paddle
             	              NSBallYAdd <= 4;
             	              NSWallVec <= "0000000000000011111" & CSWallVec(12 downto 0);      -- FIXME 
             	          end if;
             	      end if;
             	      
                   elsif CSBallYAdd <= 13 then                                                  -- against left wall
                      zone <= 5;
                      if CSBallDir(2) = '1' then
                          NSBallXAdd <= CSBallXAdd - 1;                                         -- NW -> NE 
             	          NSBallYAdd <= CSBallYAdd + 1;
             	          NsBallDir <= "101";
             	      else
             	          NSBallXAdd <= CSBallXAdd - 1;                                         -- SW -> SE
             	          NSBallYAdd <= CSBallYAdd - 1;
             	          NsBallDir <= "001";
             	      end if;
             	      
                   else                                                                         -- below top wall in left corner
                      zone <= 9;
                      NSBallXAdd <= CSBallXAdd - 1;                                             -- SE
             	      NSBallYAdd <= CSBallYAdd - 1;
             	      NsBallDir <= "001";
             	      add	<= "010" & "01111";                                                 -- reg32x32 row 15 (wall row) 
                      if reg32x32_dOut(31) = '1' then                                           -- if wall piece we increment score and remove it
                          NSScore <= CSScore + 1;
                          NSWallVec <= "0" & CSWallVec(30 downto 0);
                      end if;
                   end if;
                   
                   
               elsif CSBallXAdd = 0 then                                                        -- right wall
                   if CSBallYAdd = 4 then                                                       -- above paddle in right corner
                      zone <= 10;
                      add	<= "010" & "00010";                                                 -- paddle row
                      if reg32x32_dOut(31) = '1' then                                           -- if paddle
                          NSBallXAdd <= CSBallXAdd + 1;                                         -- NW
             	          NSBallYAdd <= CSBallYAdd + 1;
             	          NsBallDir <= "110";
             	      else                                                                      -- else we lose a life
             	          NSLives <= CSLives - 1;
             	          if NSLives > 0 then                                                   -- if we have more lives, reset ball and paddle
             	              NS <= initBall;
             	              NSBallXAdd <= 16;                                                 -- ball back to middle above paddle
             	              NSBallYAdd <= 4;
             	              NSWallVec <= CSWallVec(12 downto 0) & "1111100000000000000";      -- FIXME 
             	          end if;
             	      end if;
             	      
                   elsif CSBallYAdd <= 13 then                                                  -- against right wall
                      zone <= 4;
                      if CSBallDir(2) = '1' then
                          NSBallXAdd <= CSBallXAdd + 1;                                         -- NE -> NW 
             	          NSBallYAdd <= CSBallYAdd + 1;
             	          NsBallDir <= "110";
             	      else
             	          NSBallXAdd <= CSBallXAdd + 1;                                         -- SE -> SW
             	          NSBallYAdd <= CSBallYAdd - 1;
             	          NsBallDir <= "010";
             	      end if;
             	      
                   else                                                                         -- below top wall in right corner
                      zone <= 8;
                      NSBallXAdd <= CSBallXAdd + 1;                                             -- SW
             	      NSBallYAdd <= CSBallYAdd - 1;
             	      NsBallDir <= "010";
             	      add	<= "010" & "01111";                                                 -- reg32x32 row 15 (wall row) 
                      if reg32x32_dOut(0) = '1' then                                            -- if wall piece we increment score and remove it
                          NSScore <= CSScore + 1;
                          NSWallVec <= CSWallVec(31 downto 1) & "0";
                      end if;
                   end if;
                   

               elsif CSBallYAdd = 14 then                                                       -- just below top wall
                   zone <= 3;
                   case CSBallDir(1 downto 0) is                                                -- 00 we go straight down, 11 not valid, will not occur
                       when "01"   =>                                                           -- if NE, we bounce to SE 
                           NSBallXAdd <= CSBallXAdd - 1;                                        
                           NSBallYAdd <= CSBallYAdd - 1;
                           NsBallDir <= "001";
                       when "10"   => NSBallXAdd <= CSBallXAdd + 1;                             -- if NW, we bounce to SW 
                           NSBallXAdd <= CSBallXAdd + 1;
                           NSBallYAdd <= CSBallYAdd - 1;
                           NsBallDir <= "010";
                       when others => 
                           NSBallYAdd <= CSBallYAdd - 1;
                           NsBallDir <= "000"; 
                   end case;
                   if (CSBallVec and CSWallVec) > "0" then                                      -- if there was a wall piece infront of the ball, we remove it and increment score
                       NSScore <= CSScore + 1;
                       NSWallVec <= (CSBallVec xor CSWallVec);                                  -- since we ANDed first, we can XOR our ball and wall
                   end if;
                   
                   
               else                                                                             -- just above paddle
                   zone <= 2;
                   if (CSBallVec and CSPaddleVec) > "0" then                                    -- if paddle and ball beside each other
                       add	<= "010" & "00010";
             	       NSBallYAdd <= CSBallYAdd + 1;
             	       NsBallDir <= "100";    
                       -- TODO either shift anded signal of ball and paddle. or . add in new signal for LSBXadd of paddle
                   else                                                                         -- else we lose a lfe
                      NSLives <= CSLives - 1;
                      if NSLives > 0 then                                                       -- if we have more lifes reset ball and paddle
             	          NS <= initBall;
             	          NSBallXAdd <= 16;                                                     -- ball back to middle above paddle
             	          NSBallYAdd <= 4;
                          NSWallVec <= "00000000000000111110000000000000";                      -- FIXME 
                      end if;
                   end if;
			       
			   end if;
			   
			   if NSLives = 0 then                                                               -- if no more lives, we end game
			       NS <= endGame;
			   else                                                                              -- else write stuff to mem and loop around again
			       if NSScore > CSScore then
			           wr   	      <= '1';
			           add	          <= "010" & "00000";               -- reg32x32 row 0 
			           datToMem      <= X"000000" & "000" & std_logic_vector( to_unsigned(NSScore, 5) );
			       end if;
			       if NSLives < CSLives then
			           wr   	      <= '1';
			           add	          <= "010" & "00001";               -- reg32x32 row 1 
			           datToMem      <= X"000000" & "000" & std_logic_vector( to_unsigned(NSLives, 5) );
			       end if;                                                                              
			       NS <= writeBallToMem;
			   end if;								           
			  			   
           	else -- CSBallNumDlyCount != CSBallNumDlyMax 
	           NSBallNumDlyCount <= CSBallNumDlyCount + 1; -- increment counter
           	   NS  <= waitState;
           	end if;
 
		when NW =>                                                          -- BB State for NW Direction
             NSBallXAdd <= CSBallXAdd + 1;                                         
             NSBallYAdd <= CSBallYAdd + 1;
             NsBallDir <= "110";		
			 NS <= writeBallToMem;		
      
		when N =>                                                           -- BB State for N Direction
             NSBallXAdd <= CSBallXAdd;                                         
             NSBallYAdd <= CSBallYAdd + 1;
             NsBallDir <= "";     		
			 NS <= writeBallToMem;		
			 
		when NE =>                                                          -- BB State for NE active 
             NSBallXAdd <= CSBallXAdd - 1;                                         
             NSBallYAdd <= CSBallYAdd + 1;
             NsBallDir <= "101";                                                            
			 NS <= writeBallToMem;		
			 			 
		when SE =>                                                          -- BB State for SE Direction
             NSBallXAdd <= CSBallXAdd - 1;                                         
             NSBallYAdd <= CSBallYAdd - 1;
             NsBallDir <= "001";		
			 NS <= writeBallToMem;		
			 
		when S =>                                                           -- BB State for S Direction
             NSBallXAdd <= CSBallXAdd; 
             NSBallYAdd <= CSBallYAdd - 1;
             NsBallDir <= "";	
			 NS <= writeBallToMem;	
			 	
		when SW =>                                                          -- BB State for S Direction
             NSBallXAdd <= CSBallXAdd + 1;
             NSBallYAdd <= CSBallYAdd - 1;
             NsBallDir <= "010";		
			 NS <= writeBallToMem;				 
			 
		when writeBallToMem =>                                                           -- write new ball row
             wr                       <= '1'; 					        			      
             add(7 downto 5)          <= "010";                                          -- reg32x32 memory bank select 
             add(4 downto 0)          <= std_logic_vector( to_unsigned(CSBallYAdd, 5) ); -- row address
	   		 datToMem                 <= (others => '0');							     -- clear vector  
   	         datToMem( to_integer(to_unsigned(CSBallXAdd, 5)) ) <= '1';                  -- ball bit asserted, FIXME Why dont we write next state ball to mem?
			 NS <= writeWallToMem;
			 
	    when writeWallToMem =>         --FIXME is the best decision?                                                  -- write new Wall row
             wr   	       <= '1';
			 add           <= "010" & "01111";               -- reg32x32 row 15
			 datToMem      <= CSWallVec;
			 NS <= waitState;
		

		when endGame =>                          
			-- <perform pattern write to arena to indicate game over>
           	NS            <= writeToCSR0;            -- finish. Return done state and return control to host  TODO
  
		when others => 
			null;
	end case;
end process; 


-- Synchronous process registering current FSM state value, and other registered signals
-- registers include chip enable control
stateReg_i: process (clk, rst)
begin
  if rst = '1' then 		
    CS 	                <= idle;		
	CSWallVec           <= (others => '0');
	CSBallVec           <= (others => '0');
	CSPaddleVec         <= (others => '0');
    CSBallXAdd          <= 0;
    CSBallYAdd          <= 0;
    CSBallDir           <= (others => '0');
    CSScore             <= 0;
    CSLives             <= 0;
    CSDlyCount          <= 0;
    CSPaddleNumDlyCount <= 0;
    CSBallNumDlyCount   <= 0;
    CSDlyCountMax       <= 0;
    CSDlyCount          <= 0;
    CSPaddleNumDlyMax   <= 0;
	CSBallNumDlyMax     <= 0;
  elsif clk'event and clk = '1' then 
    if ce = '1' then
		CS 	                <= NS;		
		CSWallVec           <= NSWallVec;      
		CSBallVec           <= NSBallVec;      
		CSPaddleVec         <= NSPaddleVec;    
		CSBallXAdd          <= NSBallXAdd;     
		CSBallYAdd          <= NSBallYAdd;     
		CSBallDir           <= NSBallDir;      
		CSScore             <= NSScore;        
		CSLives             <= NSLives;        
		CSDlyCount          <= NSDlyCount;           
		CSPaddleNumDlyCount <= NSPaddleNumDlyCount;
		CSBallNumDlyCount   <= NSBallNumDlyCount; 
        CSDlyCountMax       <= NSDlyCountMax;
        CSDlyCount          <= NSDlyCount;
		CSPaddleNumDlyMax   <= NSPaddleNumDlyMax;
		CSBallNumDlyMax     <= NSBallNumDlyMax;
     end if;
  end if;
end process; 

end RTL;